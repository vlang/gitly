module highlight

fn init_d() Lang {
	return Lang{
		name:            'D'
		lang_extensions: ['d']
		line_comments:   '//'
		mline_comments:  ['/*', '*/', '/+', '+/']
		string_start:    ['"', "'"]
		color:           '#ba595e'
		keywords:        [
			'abstract',
			'alias',
			'align',
			'asm',
			'assert',
			'auto',
			'bool',
			'break',
			'byte',
			'case',
			'cast',
			'catch',
			'char',
			'class',
			'const',
			'continue',
			'dchar',
			'debug',
			'default',
			'delegate',
			'deprecated',
			'do',
			'double',
			'else',
			'enum',
			'export',
			'extern',
			'false',
			'final',
			'finally',
			'float',
			'for',
			'foreach',
			'foreach_reverse',
			'function',
			'goto',
			'if',
			'immutable',
			'import',
			'in',
			'inout',
			'int',
			'interface',
			'invariant',
			'is',
			'lazy',
			'long',
			'macro',
			'mixin',
			'module',
			'new',
			'nothrow',
			'null',
			'out',
			'override',
			'package',
			'pragma',
			'private',
			'protected',
			'public',
			'pure',
			'real',
			'ref',
			'return',
			'scope',
			'shared',
			'short',
			'static',
			'struct',
			'super',
			'switch',
			'synchronized',
			'template',
			'this',
			'throw',
			'true',
			'try',
			'typeid',
			'typeof',
			'ubyte',
			'uint',
			'ulong',
			'union',
			'unittest',
			'ushort',
			'version',
			'void',
			'wchar',
			'while',
			'with',
			'__FILE__',
			'__FILE_FULL_PATH__',
			'__MODULE__',
			'__LINE__',
			'__FUNCTION__',
			'__PRETTY_FUNCTION__',
			'__gshared',
			'__traits',
			'__vector',
			'__parameters',
		]
	}
}
