module highlight

fn init_cs() Lang {
	return Lang{
		name:            'C#'
		lang_extensions: ['cs']
		line_comments:   '//'
		mline_comments:  ['/*', '*/']
		string_start:    ['"', "'"]
		color:           '#178600'
		keywords:        [
			'abstract',
			'add',
			'alias',
			'async',
			'await',
			'base',
			'bool',
			'break',
			'by',
			'byte',
			'case',
			'catch',
			'char',
			'checked',
			'class',
			'const',
			'continue',
			'decimal',
			'default',
			'delegate',
			'do',
			'double',
			'else',
			'enum',
			'event',
			'explicit',
			'extern',
			'false',
			'finally',
			'fixed',
			'float',
			'for',
			'foreach',
			'from',
			'get',
			'goto',
			'group',
			'if',
			'implicit',
			'in',
			'int',
			'interface',
			'internal',
			'is',
			'join',
			'let',
			'lock',
			'long',
			'namespace',
			'new',
			'null',
			'object',
			'operator',
			'orderby',
			'out',
			'override',
			'params',
			'partial',
			'private',
			'protected',
			'public',
			'readonly',
			'ref',
			'remove',
			'return',
			'sbyte',
			'sealed',
			'select',
			'set',
			'short',
			'sizeof',
			'stackalloc',
			'static',
			'string',
			'struct',
			'switch',
			'this',
			'throw',
			'true',
			'try',
			'typeof',
			'uint',
			'ulong',
			'unchecked',
			'unsafe',
			'ushort',
			'using',
			'value',
			'var',
			'virtual',
			'void',
			'volatile',
			'where',
			'while',
			'yield',
		]
	}
}
