module api

pub struct ApiCommitCount {
	ApiResponse
pub:
	result int
}
