module main

const (
	ignored_folder = ['thirdparty']
)
