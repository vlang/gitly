// Copyright (c) 2019-2020 Alexander Medvednikov. All rights reserved.
// Use of this source code is governed by a GPL license that can be found in the LICENSE file.
module main

import os
import time

struct Branch {
mut:
	id     int
	repo_id int
	name   string // branch name
	author string // author of latest commit on branch
	hash   string // hash of latest commit on branch
	date   int // time of latest commit on branch
}

fn (mut app App) fetch_branches(r Repo) {
	mut branch := Branch{}
	current := os.getwd()
	os.chdir(r.git_dir)
	data := r.git('branch -a')
	for remote_branch in data.split_into_lines() {
		if remote_branch.contains('remotes/') && !remote_branch.contains('HEAD') {
			temp_branch := remote_branch.trim_space().after('remotes/')
			_ := r.git('checkout -t $temp_branch')
			branch.repo_id = r.id
			branch.name = temp_branch.after('origin/')
			hash_data := os.read_lines('.git/refs/heads/$branch.name') or {
				app.error('Error: $err')
				return
			}
			branch.hash = hash_data[0].substr(0, 7)
			branch_data := r.git('log -1 --pretty="%aE$log_field_separator%cD" $branch.hash')
			args := branch_data.split(log_field_separator)
			branch.author = args[0]
			date := time.parse_rfc2822(args[1]) or {
				app.error('Error: $err')
				return
			}
			branch.date = int(date.unix)
			app.insert_branch(branch)
		}
	}
	_ := r.git('checkout master')
	os.chdir(current)
}

fn (branch Branch) relative() string {
	return time.unix(branch.date).relative()
}

fn (mut app App) insert_branch(branch Branch) {
	sql app.db {
		insert branch into Branch
	}
}

fn (mut app App) find_branches_by_repo_id(repo_id int) []Branch {
	return sql app.db {
		select from Branch where repo_id == repo_id
	}
}

fn (mut app App) count_of_branches_by_repo_id(repo_id int) int {
	return sql app.db {
		select count from Branch where repo_id == repo_id
	}
}
