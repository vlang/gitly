module api

pub struct ApiIssueCount {
	ApiResponse
pub:
	result int
}
