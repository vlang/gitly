module api

struct ApiResponse {
pub:
	success bool
}
