// Copyright (c) 2020 Alexander Medvednikov. All rights reserved.
// Use of this source code is governed by a GPL license that can be found in the LICENSE file.
module main

import vweb
import time
import rand
import math
import libsodium
import encoding.base64

['/login']
pub fn (mut app App) login() vweb.Result {
	random_seed()
	csrf := rand.string(30)
	app.set_cookie({
		name: 'csrf'
		value: csrf
	})
	if app.logged_in() {
		return app.not_found()
	}
	return $vweb.html()
}

[post]
['/login']
pub fn (mut app App) handle_login() vweb.Result {
	if app.settings.only_gh_login {
		return app.r_home()
	}
	username := app.form['username']
	password := app.form['password']
	if username == '' || password == '' {
		return app.redirect('/login')
	}
	user := app.find_user_by_username(username) or {
		return app.redirect('/login')
	}
	if user.is_blocked {
		return app.redirect('/login')
	}
	if !check_password(password, username, user.password) {
		app.inc_user_login_attempts(user.id)
		if user.login_attempts == max_login_attempts {
			app.warn('User $user.username got blocked')
			app.block_user(user.id)
		}
		return app.redirect('/login')
	}
	if !user.is_registered {
		return app.redirect('/login')
	}
	ip := app.client_ip(user.id.str()) or {
		return app.r_home()
	}
	app.auth_user(user, ip)
	app.security_log({
		user_id: user.id
		kind: .logged_in
	})
	return app.r_home()
}

pub fn (mut app App) auth_user(user User, ip string) {
	_ := time.utc().add_days(expire_length)
	// token := if user.token == '' { app.add_token(user.id) } else { user.token }
	token := app.add_token(user.id, ip)
	println(token)
	app.update_user_login_attempts(user.id, 0)
	// println('cookie: setting token=$token id=$user.id')
	expire_date := time.now().add_days(200)
	app.set_cookie({
		name: 'id'
		value: user.id.str()
		expires: expire_date
	})
	app.set_cookie({
		name: 'token'
		value: token
		expires: expire_date
	})
	// app.set_cookie_with_expire_date('id', user.id.str(), expires)
	// app.set_cookie_with_expire_date('token', token, expires)
}

pub fn (mut app App) logged_in() bool {
	id := app.get_cookie('id') or {
		return false
	}
	token := app.get_cookie('token') or {
		return false
	}
	ip := app.client_ip(id) or {
		return false
	}
	t := app.find_user_token(id.int(), ip)
	blocked := app.check_user_blocked(id.int())
	if blocked {
		app.logout()
		return false
	}
	u := app.find_user_by_id(id.int()) or { return false }
	//de_cry := libsodium.new_secret_box(u.key).decrypt_string(base64.decode(token).bytes())
	return id != '' && token != '' && t != '' && base64.decode(token) == t /*libsodium.new_secret_box(u.key).decrypt_string(token.bytes()) == t*/
}

pub fn (mut app App) logout() vweb.Result {
	app.set_cookie({
		name: 'id'
		value: ''
	})
	app.set_cookie({
		name: 'token'
		value: ''
	})
	return app.r_home()
}

pub fn (mut app App) get_user_from_cookies() ?User {
	id := app.get_cookie('id') or {
		return none
	}
	token := app.get_cookie('token') or {
		return none
	}
	mut user := app.find_user_by_id(id.int()) or {
		return none
	}
	ip := app.client_ip(id) or {
		return none
	}
	if base64.decode(token) != app.find_user_token(user.id, ip) {
		return none
	}
	user.b_avatar = user.avatar != ''
	if !user.b_avatar {
		user.avatar = user.username.bytes()[0].str()
	}
	return user
}

['/register']
pub fn (mut app App) register() vweb.Result {
	if app.settings.only_gh_login {
		return app.r_home()
	}
	app.path = ''
	return $vweb.html()
}

[post]
['/register']
pub fn (mut app App) handle_register() vweb.Result {
	if app.settings.only_gh_login {
		return app.r_home()
	}
	username := app.form['username']
	if username in ['login', 'register', 'new', 'new_post', 'oauth'] {
		app.error('Username `$username` is not available')
		return app.register()
	}
	user_chars := username.bytes()
	if user_chars.len > max_username_len {
		app.error('Username is too long (max. $max_username_len)')
		return app.register()
	}
	if username.contains('--') {
		app.error('Username cannot contain two hyphens')
		return app.register()
	}
	if user_chars[0] == `-` || user_chars.last() == `-` {
		app.error('Username cannot begin or end with a hyphen')
		return app.register()
	}
	for char in user_chars {
		if !char.is_letter() && !char.is_digit() && char != `-` {
			app.error('Username cannot contain special characters')
			return app.register()
		}
	}
	if app.form['password'] == '' {
		app.error('Password cannot be empty')
		return app.register()
	}
	password := make_password(app.form['password'], username)
	email := app.form['email']
	if username == '' || email == '' {
		app.error('Username or Email cannot be emtpy')
		return app.register()
	}
	if !app.add_user(username, password, [email], false) {
		app.error('Failed to register')
		return app.register()
	}
	user := app.find_user_by_username(username) or {
		app.error('User already exists')
		return app.register()
	}
	println('register: logging in')
	ip := app.client_ip(user.id.str()) or {
		app.error('Failed to register')
		return app.register()
	}
	app.auth_user(user, ip)
	app.security_log({
		user_id: user.id
		kind: .registered
	})
	app.settings.only_gh_login = true
	return app.redirect('/' + username)
}

fn gen_uuid_v4ish() string {
	random_seed()
	return rand.uuid_v4()
}

fn random_seed() {
	rand.seed([u32(math.floor(math.sin(time.now().unix/2)*1000)), u32(math.floor(math.cos(time.now().unix/2)*1000))])
}
