module main

struct Release {
	tag Tag
	notes string
}
